module fifo #(
   DEPTH = 16
) (
   wishbone.device wb_in,
   wishbone.controller wb_out,
);
   
   
endmodule
