package types;

   typedef struct packed {
      logic red;
      logic green;
      logic blue;
   } rgb_led_t;


endpackage
