module debug_buttons(
   input [3:0]	       buttons, switches,
   wishbone.controller wb
);

   
   
   
   
 
endmodule
  
